module test(
	input		sysclk,
	input		sys_rst,
	output		oled
);

endmodule 

